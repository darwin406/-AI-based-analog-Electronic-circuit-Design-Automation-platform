
****curciut C****

****curciut C****
.param W1=2e-07
.param W2=1.8e-07
.param W3= 3e-06
.param W4=1.8e-07
.param W5=1.8000000000000002e-07
.param W6=1.8000000000000002e-07

.param VGS = 1


V0 power GND 2
V2 Vin2 GND dc 0.978 ac 1
V1 Vin1 GND 1

*M1 Drain Gate Source Body
M1 M1G M1G power power PMOS_MODEL l=150e-9 w=1.8000000000000002e-07
M2 M2D M1G power power PMOS_MODEL l=150e-9 w=1.8000000000000002e-07
M3 M1G Vin1 M3S M3S NMOS_MODEL l=150e-9 w=5.588325445353986e-07
M4 M2D Vin2 M3S M3S NMOS_MODEL l=150e-9 w=5.588325445353986e-07
M5 output M2D power power PMOS_MODEL l=150e-9 w=1.0885876393318177e-06
M6 M6D M6D GND GND NMOS_MODEL l=150e-9 w=1.8000000000000002e-07
M7 M3S M6D GND GND NMOS_MODEL l=150e-9 w=1.8000000000000002e-07
M8 output M6D GND GND NMOS_MODEL l=150e-9 w=1.8000000000000002e-07

R1 power M6D 20k
R2 C1R2 output 20k
C1 M2D C1R2 0.5p
C2 output GND 1p

.model NMOS_MODEL NMOS level=54 version=4.7
.model PMOS_MODEL PMOS level=54 version=4.7

***********Analysis**********
.control
****DC Analysis****
op
let power_m1 = v(power) * @M1[id]
print power_m1
wrdata simulation_log/power_data.txt power_m1


****DC Sweep *****
dc V2 0 2 0.001
plot v(output)
wrdata simulation_log/dc_sweep_data.txt v(output)



* *****AC / Frequency response ****
ac dec 100 1 100G
plot vdb(output) 
print vdb(output)[0]
plot ph(output)*180/pi
wrdata simulation_log/ac_analysis_data.txt vdb(output) ph(output)

.endc
.end
    